CLK_IN_inst : CLK_IN PORT MAP (
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
